* D:\workspace\PriorityEncoder\PriorityEncoder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/01/21 12:25:11

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  GND Net-_U2-Pad2_ GND GND Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ GND Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ adc_bridge_8		
v1  Net-_U2-Pad2_ GND DC		
v2  Net-_U2-Pad5_ GND DC		
v3  Net-_U2-Pad6_ GND DC		
v4  Net-_U2-Pad7_ GND DC		
R3  Net-_R3-Pad1_ GND 1K		
R2  Net-_R2-Pad1_ GND 1K		
R1  Net-_R1-Pad1_ GND 1K		
U4  Net-_R1-Pad1_ plot_v1		
U5  Net-_R2-Pad1_ plot_v1		
U6  Net-_R3-Pad1_ plot_v1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ PriorityEncoder		
U3  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_R3-Pad1_ Net-_R2-Pad1_ Net-_R1-Pad1_ dac_bridge_3		

.end
